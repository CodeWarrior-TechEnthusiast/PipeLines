`include "define.v"

module EXE_WB_stage (
	
	input  clk,  rst,
	
);




//EXE_WWB register to save the values.


endmodule


