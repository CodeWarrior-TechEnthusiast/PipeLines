`include "define.v"

module ID_EXE_stage (
	
	input  clk,  rst, 

	
);



//Here we need not take write enable (wen) as it is always 1 for R and I type instructions.
//ID_EXE register to save the values.



endmodule


