`timescale 1ns / 1ps
`include "define.v"

module pipelined_3stage(clk, rst, aluout);

input clk;				
											
input rst;

output [`DSIZE-1:0] aluout;	

 
endmodule


