`timescale 1ns / 1ps
`include "define.v"

module pipelined_regfile_4stage(clk, rst, aluout_EXE_WB);

input clk;				
											
input	rst;

	
output [`DSIZE-1:0] aluout_EXE_WB;								
 	 


endmodule


